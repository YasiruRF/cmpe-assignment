library verilog;
use verilog.vl_types.all;
entity MainALU_vlg_vec_tst is
end MainALU_vlg_vec_tst;
