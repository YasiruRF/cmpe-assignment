library verilog;
use verilog.vl_types.all;
entity RightShift_vlg_vec_tst is
end RightShift_vlg_vec_tst;
