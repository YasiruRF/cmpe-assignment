library verilog;
use verilog.vl_types.all;
entity AndOrXorXnor_vlg_vec_tst is
end AndOrXorXnor_vlg_vec_tst;
