library verilog;
use verilog.vl_types.all;
entity fourbitAU_vlg_vec_tst is
end fourbitAU_vlg_vec_tst;
