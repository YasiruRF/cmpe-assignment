library verilog;
use verilog.vl_types.all;
entity AmultiplyB_vlg_vec_tst is
end AmultiplyB_vlg_vec_tst;
