library verilog;
use verilog.vl_types.all;
entity RotateRight_vlg_vec_tst is
end RotateRight_vlg_vec_tst;
