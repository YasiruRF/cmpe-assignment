library verilog;
use verilog.vl_types.all;
entity LeftShift_vlg_vec_tst is
end LeftShift_vlg_vec_tst;
