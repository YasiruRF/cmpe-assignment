library verilog;
use verilog.vl_types.all;
entity RotateLeft_vlg_vec_tst is
end RotateLeft_vlg_vec_tst;
