library verilog;
use verilog.vl_types.all;
entity LogicalUnitMain_vlg_vec_tst is
end LogicalUnitMain_vlg_vec_tst;
