library verilog;
use verilog.vl_types.all;
entity Transfer_vlg_vec_tst is
end Transfer_vlg_vec_tst;
