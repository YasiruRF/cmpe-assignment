library verilog;
use verilog.vl_types.all;
entity ArithmaticRightShift_vlg_vec_tst is
end ArithmaticRightShift_vlg_vec_tst;
